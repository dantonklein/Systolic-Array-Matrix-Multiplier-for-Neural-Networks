module controller (
    
);


endmodule